module vimgui

